module lab5(num2, num1, num0);
	output [6:0] num2, num1, num0;
	
	assign num2 = 7'b1111001; //1
	assign num1 = 7'b1111001; //1
	assign num0 = 7'b1111000; //7
	
endmodule
